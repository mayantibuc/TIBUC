CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 110 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
76546066 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 83 180 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6986 0 0
2
5.89883e-315 0
0
9 CC 7-Seg~
183 1023 161 0 9 19
10 17 16 15 14 13 12 11 18 19
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
8745 0 0
2
5.89883e-315 0
0
7 Pulser~
4 166 343 0 10 12
0 20 21 9 22 0 0 5 5 2
7
0
0 0 4640 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9592 0 0
2
5.89883e-315 5.26354e-315
0
9 2-In AND~
219 588 80 0 3 22
0 3 5 7
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
8748 0 0
2
5.89883e-315 5.30499e-315
0
9 2-In AND~
219 453 70 0 3 22
0 2 4 3
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7168 0 0
2
5.89883e-315 5.32571e-315
0
2 +V
167 164 112 0 1 3
0 10
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
631 0 0
2
5.89883e-315 5.34643e-315
0
6 74LS48
188 837 201 0 14 29
0 6 5 4 2 23 24 11 12 13
14 15 16 17 25
0
0 0 4832 0
7 74LS248
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9466 0 0
2
5.89883e-315 5.36716e-315
0
6 74112~
219 655 215 0 7 32
0 10 7 9 7 10 26 6
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
3266 0 0
2
5.89883e-315 5.37752e-315
0
6 74112~
219 514 217 0 7 32
0 10 3 9 3 10 27 5
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
7693 0 0
2
5.89883e-315 5.38788e-315
0
6 74112~
219 377 218 0 7 32
0 10 2 9 2 10 28 4
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U1B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
3723 0 0
2
5.89883e-315 5.39306e-315
0
6 74112~
219 244 214 0 7 32
0 10 8 9 8 10 29 2
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
3440 0 0
2
5.89883e-315 5.39824e-315
0
37
1 0 2 0 0 8192 0 5 0 0 14 3
429 61
335 61
335 182
0 4 2 0 0 0 0 0 10 14 0 3
318 180
318 200
353 200
3 4 3 0 0 4224 0 5 9 0 0 3
474 70
474 199
490 199
0 3 4 0 0 8320 0 0 7 13 0 5
415 180
415 300
749 300
749 183
805 183
4 0 2 0 0 12416 0 7 0 0 14 5
805 192
761 192
761 135
307 135
307 180
2 0 5 0 0 12416 0 7 0 0 10 5
805 174
732 174
732 285
555 285
555 181
7 1 6 0 0 12416 0 8 7 0 0 4
679 179
729 179
729 165
805 165
0 4 7 0 0 8192 0 0 8 9 0 3
609 179
609 197
631 197
3 2 7 0 0 4224 0 4 8 0 0 3
609 80
609 179
631 179
7 2 5 0 0 0 0 9 4 0 0 4
538 181
555 181
555 89
564 89
2 0 3 0 0 0 0 9 0 0 12 3
490 181
481 181
481 70
1 3 3 0 0 0 0 4 5 0 0 3
564 71
564 70
474 70
7 2 4 0 0 0 0 10 5 0 0 4
401 182
415 182
415 79
429 79
7 2 2 0 0 0 0 11 10 0 0 6
268 178
307 178
307 180
318 180
318 182
353 182
4 0 8 0 0 4224 0 11 0 0 16 3
220 196
150 196
150 180
2 1 8 0 0 0 0 11 1 0 0 4
220 178
150 178
150 180
95 180
3 0 9 0 0 4096 0 11 0 0 21 2
214 187
214 334
3 0 9 0 0 0 0 10 0 0 21 4
347 191
347 319
349 319
349 334
3 0 9 0 0 0 0 9 0 0 21 4
484 190
484 319
485 319
485 334
3 0 9 0 0 0 0 8 0 0 21 4
625 188
625 319
619 319
619 334
3 0 9 0 0 4224 0 3 0 0 0 2
190 334
733 334
5 0 10 0 0 4096 0 11 0 0 30 2
244 226
244 259
5 0 10 0 0 0 0 10 0 0 30 4
377 230
377 244
379 244
379 259
5 0 10 0 0 0 0 9 0 0 30 4
514 229
514 244
515 244
515 259
5 0 10 0 0 0 0 8 0 0 30 4
655 227
655 244
649 244
649 259
1 0 10 0 0 0 0 8 0 0 30 4
655 152
655 136
649 136
649 121
1 0 10 0 0 0 0 9 0 0 30 4
514 154
514 136
515 136
515 121
1 0 10 0 0 0 0 10 0 0 30 4
377 155
377 136
379 136
379 121
1 0 10 0 0 0 0 11 0 0 30 2
244 151
244 121
1 0 10 0 0 12416 0 6 0 0 0 4
164 121
719 121
719 259
141 259
7 7 11 0 0 12416 0 2 7 0 0 6
1038 197
1037 197
1037 269
904 269
904 165
869 165
6 8 12 0 0 12416 0 2 7 0 0 6
1032 197
1031 197
1031 259
918 259
918 174
869 174
5 9 13 0 0 12416 0 2 7 0 0 6
1026 197
1025 197
1025 251
925 251
925 183
869 183
4 10 14 0 0 20608 0 2 7 0 0 6
1020 197
1019 197
1019 243
945 243
945 192
869 192
3 11 15 0 0 20608 0 2 7 0 0 6
1014 197
1013 197
1013 232
968 232
968 201
869 201
2 12 16 0 0 20608 0 2 7 0 0 6
1008 197
1007 197
1007 226
979 226
979 210
869 210
13 1 17 0 0 4224 0 7 2 0 0 4
869 219
1001 219
1001 197
1002 197
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
268 403 415 425
277 410 405 426
16 Tibuc, May An M.
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
